megawizard_vjtag_inst : megawizard_vjtag PORT MAP (
		ir_out	 => ir_out_sig,
		tdo	 => tdo_sig,
		ir_in	 => ir_in_sig,
		tck	 => tck_sig,
		tdi	 => tdi_sig,
		virtual_state_cdr	 => virtual_state_cdr_sig,
		virtual_state_cir	 => virtual_state_cir_sig,
		virtual_state_e1dr	 => virtual_state_e1dr_sig,
		virtual_state_e2dr	 => virtual_state_e2dr_sig,
		virtual_state_pdr	 => virtual_state_pdr_sig,
		virtual_state_sdr	 => virtual_state_sdr_sig,
		virtual_state_udr	 => virtual_state_udr_sig,
		virtual_state_uir	 => virtual_state_uir_sig
	);
